module hex16seg (hex, display);
	input [15:0] hex;
	output [0:15] display;

	reg [0:15] display;

	/*
	 *       0  
	 *      ---  
	 *     |   |
	 *    5|   |1
	 *     | 6 |
	 *      ---  
	 *     |   |
	 *    4|   |2
	 *     |   |
	 *      ---  
	 *       3  
	 */
	always @ (hex)
		case (hex)
			16'b000000000000000: display = 16'b0000000000000001; //0
			16'b000000000000001: display = 16'b0000000001001111; //1
			16'b000000000000010: display = 16'b0000000000010010; //2
			16'b000000000000011: display = 16'b0000000000000110; //3
			16'b000000000000100: display = 16'b0000000001001100; //4
			16'b000000000000101: display = 16'b0000000000100100; //5
			16'b000000000000110: display = 16'b0000000000100000; //6
			16'b000000000000111: display = 16'b0000000000001111; //7
			16'b000000000001000: display = 16'b0000000000000000; //8
			16'b000000000001001: display = 16'b0000000000000100; //9
			16'b000000000001010: display = 16'b0000000000001000; //A
			16'b000000000001011: display = 16'b0000000001100000; //B
			16'b000000000001100: display = 16'b0000000000110001; //C
			16'b000000000001101: display = 16'b0000000001000010; //D
			16'b000000000001110: display = 16'b0000000000110000; //E
			16'b000000000001111: display = 16'b0000000000111000; //F
		endcase
endmodule